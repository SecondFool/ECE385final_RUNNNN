module player1(input [9:0] pX,
				input [9:0] pY,
				input [31:0] f1,
				output logic [2:0] cidx
				);
			
	
	//logic [2:0] IMG [899:0] = '{3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b010,3'b011,3'b010,3'b010,3'b010,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b011,3'b011,3'b010,3'b100,3'b100,3'b100,3'b100,3'b011,3'b100,3'b100,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b011,3'b010,3'b010,3'b010,3'b011,3'b011,3'b010,3'b100,3'b100,3'b011,3'b011,3'b011,3'b100,3'b100,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b011,3'b011,3'b010,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b011,3'b010,3'b011,3'b010,3'b010,3'b011,3'b010,3'b100,3'b010,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b100,3'b011,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b011,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b011,3'b010,3'b010,3'b011,3'b011,3'b011,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b011,3'b010,3'b011,3'b011,3'b011,3'b011,3'b100,3'b000,3'b011,3'b011,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b101,3'b000,3'b000,3'b000,3'b000,3'b011,3'b011,3'b011,3'b011,3'b011,3'b100,3'b100,3'b100,3'b011,3'b011,3'b011,3'b010,3'b010,3'b010,3'b011,3'b100,3'b100,3'b011,3'b010,3'b100,3'b010,3'b010,3'b000,3'b101,3'b101,3'b101,3'b101,3'b110,3'b110,3'b000,3'b011,3'b011,3'b011,3'b011,3'b011,3'b100,3'b001,3'b100,3'b100,3'b100,3'b010,3'b010,3'b011,3'b001,3'b100,3'b100,3'b010,3'b100,3'b010,3'b010,3'b010,3'b010,3'b000,3'b101,3'b101,3'b101,3'b110,3'b110,3'b110,3'b110,3'b000,3'b000,3'b011,3'b011,3'b011,3'b100,3'b001,3'b100,3'b011,3'b011,3'b010,3'b001,3'b001,3'b011,3'b011,3'b010,3'b010,3'b010,3'b100,3'b100,3'b010,3'b010,3'b000,3'b101,3'b101,3'b101,3'b110,3'b101,3'b110,3'b110,3'b110,3'b000,3'b011,3'b011,3'b011,3'b011,3'b001,3'b100,3'b011,3'b100,3'b010,3'b001,3'b011,3'b010,3'b010,3'b010,3'b100,3'b010,3'b100,3'b010,3'b010,3'b010,3'b000,3'b101,3'b101,3'b101,3'b110,3'b101,3'b110,3'b110,3'b110,3'b110,3'b000,3'b011,3'b011,3'b011,3'b011,3'b010,3'b010,3'b010,3'b011,3'b011,3'b011,3'b011,3'b010,3'b100,3'b010,3'b010,3'b100,3'b010,3'b010,3'b010,3'b000,3'b101,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b011,3'b011,3'b011,3'b011,3'b011,3'b011,3'b011,3'b011,3'b010,3'b010,3'b100,3'b010,3'b010,3'b100,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b101,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b011,3'b010,3'b011,3'b011,3'b010,3'b010,3'b011,3'b001,3'b100,3'b100,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b101,3'b101,3'b110,3'b110,3'b101,3'b110,3'b110,3'b110,3'b110,3'b011,3'b011,3'b011,3'b011,3'b011,3'b100,3'b100,3'b001,3'b001,3'b100,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b101,3'b101,3'b101,3'b110,3'b101,3'b110,3'b110,3'b110,3'b011,3'b011,3'b011,3'b010,3'b011,3'b011,3'b011,3'b001,3'b011,3'b011,3'b010,3'b001,3'b011,3'b010,3'b100,3'b100,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b101,3'b101,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b011,3'b011,3'b011,3'b011,3'b011,3'b011,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b011,3'b010,3'b100,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b101,3'b101,3'b101,3'b101,3'b110,3'b110,3'b110,3'b000,3'b011,3'b011,3'b011,3'b011,3'b011,3'b100,3'b011,3'b100,3'b100,3'b100,3'b010,3'b010,3'b011,3'b011,3'b100,3'b100,3'b010,3'b100,3'b100,3'b010,3'b010,3'b000,3'b000,3'b101,3'b101,3'b101,3'b000,3'b000,3'b000,3'b000,3'b011,3'b011,3'b010,3'b010,3'b010,3'b100,3'b100,3'b100,3'b011,3'b011,3'b010,3'b010,3'b001,3'b011,3'b010,3'b100,3'b100,3'b100,3'b011,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b011,3'b011,3'b011,3'b010,3'b011,3'b100,3'b100,3'b011,3'b100,3'b011,3'b011,3'b010,3'b010,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b011,3'b011,3'b010,3'b011,3'b010,3'b010,3'b011,3'b011,3'b011,3'b011,3'b000,3'b000,3'b011,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b100,3'b010,3'b011,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b011,3'b010,3'b011,3'b011,3'b011,3'b011,3'b011,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b010,3'b011,3'b011,3'b011,3'b011,3'b010,3'b011,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b011,3'b011,3'b010,3'b011,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b011,3'b011,3'b011,3'b100,3'b100,3'b011,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b011,3'b010,3'b010,3'b010,3'b010,3'b010,3'b100,3'b100,3'b100,3'b011,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001};	
	logic [2:0] IMG1 [899:0] = '{3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001};
	logic [2:0] IMG2 [899:0] = '{3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b011,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b011,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b011,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b011,3'b000,3'b010,3'b000,3'b011,3'b011,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b010,3'b010,3'b000,3'b011,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001};
	logic [2:0] IMG3 [899:0] = '{3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b100,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b100,3'b100,3'b100,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b010,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b100,3'b100,3'b100,3'b100,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b100,3'b100,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b000,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001};
	logic [9:0] idx;
	assign idx = pX*30 + pY;
	always_comb
		begin
			case(f1)
					0:
						begin
							cidx = IMG1[899-idx];
						end
					1:
						begin
							cidx = IMG2[899-idx];
						end
					2:
						begin
							cidx = IMG3[899-idx];
						end
					3:
						begin
							cidx = IMG2[899-idx];
						end
					default:
						begin
							cidx = 0;
						end
				endcase
		end
endmodule

module player2(input [9:0] pX,
				input [9:0] pY,
				input [31:0] f2,
				output logic [2:0] cidx
				);
			
	
	logic [2:0] IMG1 [899:0] = '{3'b110,3'b000,3'b000,3'b110,3'b110,3'b000,3'b011,3'b011,3'b011,3'b011,3'b011,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b110,3'b000,3'b000,3'b110,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b011,3'b011,3'b001,3'b001,3'b011,3'b011,3'b011,3'b000,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b110,3'b110,3'b110,3'b000,3'b110,3'b110,3'b000,3'b000,3'b011,3'b011,3'b001,3'b001,3'b001,3'b011,3'b011,3'b011,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b000,3'b110,3'b110,3'b000,3'b000,3'b110,3'b000,3'b000,3'b011,3'b011,3'b011,3'b001,3'b001,3'b001,3'b011,3'b011,3'b011,3'b000,3'b000,3'b000,3'b010,3'b000,3'b010,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b110,3'b000,3'b000,3'b011,3'b011,3'b011,3'b011,3'b001,3'b001,3'b001,3'b011,3'b011,3'b000,3'b000,3'b010,3'b010,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b110,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b100,3'b100,3'b101,3'b011,3'b011,3'b011,3'b001,3'b011,3'b011,3'b011,3'b000,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b110,3'b110,3'b000,3'b000,3'b110,3'b000,3'b100,3'b100,3'b100,3'b101,3'b011,3'b011,3'b011,3'b011,3'b011,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b100,3'b101,3'b011,3'b011,3'b011,3'b101,3'b101,3'b100,3'b101,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b110,3'b000,3'b000,3'b100,3'b100,3'b100,3'b110,3'b110,3'b000,3'b000,3'b101,3'b101,3'b100,3'b110,3'b100,3'b101,3'b011,3'b100,3'b100,3'b101,3'b101,3'b100,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b100,3'b100,3'b000,3'b000,3'b101,3'b101,3'b100,3'b101,3'b000,3'b100,3'b000,3'b100,3'b101,3'b101,3'b100,3'b100,3'b101,3'b101,3'b100,3'b100,3'b101,3'b101,3'b100,3'b000,3'b101,3'b100,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b100,3'b101,3'b101,3'b001,3'b001,3'b000,3'b100,3'b100,3'b000,3'b100,3'b100,3'b100,3'b101,3'b100,3'b100,3'b101,3'b110,3'b100,3'b100,3'b101,3'b100,3'b101,3'b101,3'b100,3'b100,3'b000,3'b000,3'b000,3'b100,3'b100,3'b101,3'b101,3'b001,3'b001,3'b001,3'b101,3'b101,3'b100,3'b100,3'b000,3'b101,3'b000,3'b101,3'b100,3'b101,3'b000,3'b100,3'b100,3'b100,3'b100,3'b101,3'b110,3'b000,3'b000,3'b000,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b100,3'b001,3'b001,3'b001,3'b101,3'b101,3'b101,3'b100,3'b000,3'b101,3'b101,3'b110,3'b100,3'b100,3'b000,3'b000,3'b100,3'b000,3'b000,3'b000,3'b100,3'b101,3'b100,3'b100,3'b100,3'b100,3'b000,3'b100,3'b101,3'b101,3'b100,3'b001,3'b001,3'b101,3'b101,3'b001,3'b000,3'b100,3'b100,3'b100,3'b101,3'b110,3'b100,3'b101,3'b100,3'b000,3'b000,3'b101,3'b100,3'b101,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b101,3'b101,3'b101,3'b101,3'b101,3'b101,3'b001,3'b001,3'b000,3'b000,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b100,3'b101,3'b100,3'b100,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b101,3'b101,3'b101,3'b101,3'b101,3'b001,3'b001,3'b000,3'b000,3'b101,3'b101,3'b100,3'b101,3'b100,3'b110,3'b100,3'b101,3'b100,3'b001,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b101,3'b101,3'b101,3'b101,3'b101,3'b001,3'b001,3'b000,3'b000,3'b101,3'b100,3'b100,3'b100,3'b000,3'b100,3'b100,3'b100,3'b101,3'b001,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b101,3'b100,3'b001,3'b001,3'b101,3'b101,3'b001,3'b000,3'b100,3'b100,3'b100,3'b100,3'b101,3'b100,3'b100,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b101,3'b101,3'b100,3'b001,3'b001,3'b100,3'b101,3'b101,3'b100,3'b100,3'b100,3'b101,3'b100,3'b000,3'b100,3'b100,3'b001,3'b100,3'b001,3'b100,3'b100,3'b101,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b101,3'b001,3'b001,3'b001,3'b101,3'b101,3'b101,3'b100,3'b000,3'b100,3'b100,3'b000,3'b101,3'b100,3'b101,3'b100,3'b000,3'b101,3'b101,3'b100,3'b101,3'b100,3'b101,3'b000,3'b100,3'b100,3'b000,3'b100,3'b000,3'b100,3'b101,3'b100,3'b001,3'b001,3'b101,3'b101,3'b001,3'b000,3'b100,3'b100,3'b100,3'b100,3'b101,3'b000,3'b100,3'b000,3'b000,3'b100,3'b100,3'b101,3'b101,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b100,3'b100,3'b101,3'b101,3'b101,3'b101,3'b100,3'b000,3'b000,3'b101,3'b100,3'b101,3'b101,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b101,3'b100,3'b100,3'b100,3'b000,3'b100,3'b000,3'b100,3'b000,3'b000,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b000,3'b000,3'b100,3'b000,3'b110,3'b010,3'b010,3'b111,3'b111,3'b111,3'b111,3'b111,3'b010,3'b010,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b000,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b101,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b101,3'b111,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b110,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b101,3'b101,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b011,3'b101,3'b111,3'b010,3'b010,3'b000,3'b000,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b110,3'b000,3'b110,3'b100,3'b101,3'b100,3'b110,3'b010,3'b111,3'b111,3'b011,3'b011,3'b011,3'b011,3'b011,3'b111,3'b111,3'b010,3'b110,3'b110,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b101,3'b100,3'b101,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b011,3'b101,3'b111,3'b010,3'b010,3'b000,3'b000,3'b110,3'b110,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b101,3'b101,3'b100,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b101,3'b111,3'b111,3'b010,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b110,3'b101,3'b110,3'b010,3'b010,3'b111,3'b111,3'b111,3'b111,3'b111,3'b010,3'b000,3'b110,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b000};	
	logic [2:0] IMG2 [899:0] = '{3'b110,3'b000,3'b000,3'b110,3'b110,3'b000,3'b011,3'b011,3'b011,3'b011,3'b011,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b110,3'b000,3'b000,3'b110,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b011,3'b011,3'b001,3'b001,3'b011,3'b011,3'b011,3'b000,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b110,3'b110,3'b110,3'b000,3'b110,3'b110,3'b000,3'b000,3'b011,3'b011,3'b001,3'b001,3'b001,3'b011,3'b011,3'b011,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b000,3'b110,3'b110,3'b000,3'b000,3'b110,3'b000,3'b000,3'b011,3'b011,3'b011,3'b001,3'b001,3'b001,3'b011,3'b011,3'b011,3'b000,3'b000,3'b000,3'b010,3'b000,3'b010,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b110,3'b000,3'b000,3'b011,3'b011,3'b011,3'b011,3'b001,3'b001,3'b001,3'b011,3'b011,3'b000,3'b000,3'b010,3'b010,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b110,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b100,3'b100,3'b101,3'b011,3'b011,3'b011,3'b001,3'b011,3'b011,3'b011,3'b000,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b110,3'b110,3'b000,3'b000,3'b110,3'b000,3'b100,3'b100,3'b100,3'b101,3'b011,3'b011,3'b011,3'b011,3'b011,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b100,3'b101,3'b011,3'b011,3'b011,3'b101,3'b101,3'b100,3'b101,3'b100,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b110,3'b000,3'b000,3'b100,3'b100,3'b100,3'b110,3'b110,3'b000,3'b000,3'b101,3'b101,3'b100,3'b110,3'b100,3'b101,3'b011,3'b100,3'b100,3'b101,3'b101,3'b100,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b100,3'b100,3'b000,3'b000,3'b101,3'b101,3'b100,3'b101,3'b000,3'b100,3'b000,3'b100,3'b101,3'b101,3'b100,3'b100,3'b101,3'b101,3'b100,3'b100,3'b101,3'b101,3'b100,3'b000,3'b101,3'b100,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b000,3'b100,3'b101,3'b101,3'b001,3'b001,3'b000,3'b100,3'b100,3'b000,3'b100,3'b100,3'b100,3'b101,3'b100,3'b100,3'b101,3'b110,3'b100,3'b100,3'b101,3'b100,3'b101,3'b101,3'b100,3'b100,3'b000,3'b000,3'b000,3'b100,3'b100,3'b101,3'b101,3'b001,3'b001,3'b001,3'b101,3'b101,3'b100,3'b100,3'b000,3'b101,3'b000,3'b101,3'b100,3'b101,3'b000,3'b100,3'b100,3'b100,3'b100,3'b101,3'b110,3'b000,3'b000,3'b000,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b100,3'b001,3'b001,3'b001,3'b101,3'b101,3'b101,3'b100,3'b000,3'b101,3'b101,3'b110,3'b100,3'b100,3'b000,3'b000,3'b100,3'b000,3'b000,3'b000,3'b100,3'b101,3'b100,3'b100,3'b100,3'b100,3'b000,3'b100,3'b101,3'b101,3'b100,3'b001,3'b001,3'b101,3'b101,3'b001,3'b000,3'b100,3'b100,3'b100,3'b101,3'b110,3'b100,3'b101,3'b100,3'b000,3'b000,3'b101,3'b100,3'b101,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b101,3'b101,3'b101,3'b101,3'b101,3'b101,3'b001,3'b001,3'b000,3'b000,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b100,3'b101,3'b100,3'b100,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b101,3'b101,3'b101,3'b101,3'b101,3'b001,3'b001,3'b000,3'b000,3'b101,3'b101,3'b100,3'b101,3'b100,3'b110,3'b100,3'b101,3'b100,3'b001,3'b101,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b101,3'b101,3'b101,3'b101,3'b101,3'b001,3'b001,3'b000,3'b000,3'b101,3'b100,3'b100,3'b100,3'b000,3'b100,3'b100,3'b100,3'b101,3'b001,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b101,3'b100,3'b001,3'b001,3'b101,3'b101,3'b001,3'b000,3'b100,3'b100,3'b100,3'b100,3'b101,3'b100,3'b100,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b101,3'b101,3'b100,3'b001,3'b001,3'b100,3'b101,3'b101,3'b100,3'b100,3'b100,3'b101,3'b100,3'b000,3'b100,3'b100,3'b001,3'b100,3'b001,3'b100,3'b100,3'b101,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b101,3'b001,3'b001,3'b001,3'b101,3'b101,3'b101,3'b100,3'b000,3'b100,3'b100,3'b000,3'b101,3'b100,3'b101,3'b100,3'b000,3'b101,3'b101,3'b100,3'b101,3'b100,3'b101,3'b000,3'b100,3'b100,3'b000,3'b100,3'b000,3'b100,3'b101,3'b100,3'b001,3'b001,3'b101,3'b101,3'b001,3'b000,3'b100,3'b100,3'b100,3'b100,3'b101,3'b000,3'b100,3'b000,3'b000,3'b100,3'b100,3'b101,3'b101,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b100,3'b100,3'b101,3'b101,3'b101,3'b101,3'b100,3'b000,3'b000,3'b101,3'b100,3'b101,3'b101,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b101,3'b100,3'b100,3'b100,3'b000,3'b100,3'b000,3'b100,3'b000,3'b000,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b000,3'b000,3'b100,3'b000,3'b110,3'b010,3'b010,3'b111,3'b111,3'b111,3'b111,3'b111,3'b010,3'b010,3'b000,3'b000,3'b100,3'b100,3'b100,3'b000,3'b000,3'b100,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b101,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b101,3'b111,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b100,3'b100,3'b110,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b101,3'b101,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b011,3'b101,3'b111,3'b010,3'b010,3'b000,3'b000,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b110,3'b000,3'b110,3'b110,3'b000,3'b110,3'b100,3'b101,3'b100,3'b110,3'b010,3'b111,3'b111,3'b011,3'b011,3'b011,3'b011,3'b011,3'b111,3'b111,3'b010,3'b110,3'b110,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b101,3'b100,3'b101,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b011,3'b101,3'b111,3'b010,3'b010,3'b000,3'b000,3'b110,3'b110,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b101,3'b101,3'b100,3'b110,3'b010,3'b111,3'b111,3'b101,3'b011,3'b011,3'b101,3'b111,3'b111,3'b010,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b000,3'b000,3'b000,3'b110,3'b110,3'b101,3'b110,3'b010,3'b010,3'b111,3'b111,3'b111,3'b111,3'b111,3'b010,3'b000,3'b110,3'b000,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b000,3'b110,3'b000,3'b110,3'b000,3'b000,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b110,3'b000,3'b000,3'b000,3'b000,3'b000};	

	logic [9:0] idx;
	assign idx = pX*30 + pY;
		always_comb
		begin
			case(f2)
					0:
						begin
							cidx = IMG1[899-idx];
						end
					1:
						begin
							cidx = IMG2[899-idx];
						end
					default:
						begin
							cidx = 0;
						end
			endcase
		end
endmodule

module isplayer(input [9:0] pX,
				input [9:0] pY,
				input [9:0] pX2,
				input [9:0] pY2,
				input [9:0] DrawX,
				input [9:0] DrawY,
				output logic isp1,
				output logic isp2
	);
	always_comb
		begin
			if ((DrawX >= pX)&&(DrawX < pX+30)&&(DrawY >= pY)&&(DrawY < pY+30))
				begin
					isp1 = 1;
				end
			else
				begin
					isp1 = 0;
				end
			if ((DrawX >= pX2)&&(DrawX < pX2+30)&&(DrawY >= pY2)&&(DrawY < pY2+30))
				begin
					isp2 = 1;
				end
			else
				begin
					isp2 = 0;
				end
		end
endmodule
	
