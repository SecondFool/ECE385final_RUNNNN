module wall(input [9:0] wallX,
				input [9:0] wallY,
				input [7:0] p1ab,
				input logic isDoor,
				output logic [2:0] cidx
				);
			
	
	logic [2:0] IMG [899:0] = '{3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b010,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b001,3'b000,3'b000,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b010,3'b000,3'b001,3'b010,3'b000,3'b001,3'b000,3'b000,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b010,3'b001,3'b010,3'b000,3'b010,3'b010,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b010,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b010,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b001,3'b010,3'b001,3'b010,3'b001,3'b001,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b010,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b010,3'b010,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b010,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010};	
	logic	DOOR[899:0] = '{0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic [9:0] idx;
	assign idx = wallX*30 + wallY;
	always_comb
		begin
			if (p1ab == 1 && isDoor == 1 && DOOR[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
			else
				begin
					cidx = IMG[899 - idx];
				end
		end
endmodule


module road(input [9:0] roadX,
				input [9:0] roadY,
				input [7:0] p1ab,
				input [7:0] p2ab,
				input [1:0] SD,
				output logic [2:0] cidx
				);
			
	
	logic [2:0] IMG1 [899:0] = '{3'b100,3'b101,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b101,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b101,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b101,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b101,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b101,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b101,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b101,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b101,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b101,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b101,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b101,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b101,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b101,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100};	
	logic SHIT[899:0] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic PLANES[899:0] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic PLANED[899:0] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic [9:0] idx;
	assign idx = roadX*30 + roadY;
		always_comb
		begin
			cidx = IMG1[899 - idx];
			if (p1ab == 0 && SD == 2 && PLANES[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
			else if (p1ab == 0 && SD == 3 && PLANED[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
			else if (p2ab == 1 && SD == 1 && SHIT[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
		end
endmodule
